// Hello world in Verilog

module main;
  initial 
    begin
	
      $display("Hello, World");  //Displaying the text
      
	  $finish ;
    
	end
endmodule